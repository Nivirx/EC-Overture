module ALU (clk, rst, Instruction, A, B, D_OUT_EN, D, CF, C);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  input  wire [7:0] Instruction;
  input  wire [7:0] A;
  input  wire [7:0] B;
  output  wire [0:0] D_OUT_EN;
  output  wire [7:0] D;
  output  wire [0:0] CF;
  output  wire [7:0] C;

  TC_Splitter8 # (.UUID(64'd1753460274403159300 ^ UUID)) Splitter8_0 (.in(wire_29), .out0(wire_7), .out1(wire_82), .out2(wire_55), .out3(wire_69), .out4(wire_42), .out5(wire_31), .out6(), .out7());
  TC_Decoder3 # (.UUID(64'd812012822489249482 ^ UUID)) Decoder3_1 (.dis(1'd0), .sel0(wire_7), .sel1(wire_82), .sel2(wire_55), .out0(wire_5), .out1(wire_1), .out2(wire_4), .out3(wire_16), .out4(wire_24), .out5(wire_0), .out6(wire_26), .out7(wire_48));
  TC_Add # (.UUID(64'd1656672475853897358 ^ UUID), .BIT_WIDTH(64'd8)) Add8_2 (.in0(wire_86), .in1(wire_45), .ci(1'd0), .out(wire_33), .co(wire_21));
  TC_Switch # (.UUID(64'd2854607076807969927 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_3 (.en(wire_24), .in(wire_2), .out(wire_72));
  TC_Switch # (.UUID(64'd1098925891083976806 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_4 (.en(wire_24), .in(wire_6), .out(wire_84));
  TC_Switch # (.UUID(64'd272865694635219578 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_5 (.en(wire_24), .in(wire_62), .out(wire_22_4));
  TC_Neg # (.UUID(64'd4234413084985973774 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_6 (.in(wire_68), .out(wire_45));
  TC_Add # (.UUID(64'd2365866274018282956 ^ UUID), .BIT_WIDTH(64'd8)) Add8_7 (.in0(wire_84), .in1(wire_72), .ci(1'd0), .out(wire_62), .co(wire_23));
  TC_Switch # (.UUID(64'd2540442194520213284 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_8 (.en(wire_16), .in(wire_6), .out(wire_86));
  TC_Switch # (.UUID(64'd927777902762540353 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_9 (.en(wire_16), .in(wire_2), .out(wire_68));
  TC_Switch # (.UUID(64'd4324181735425917878 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_10 (.en(wire_16), .in(wire_33), .out(wire_22_2));
  TC_Switch # (.UUID(64'd1224106639434152846 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_11 (.en(wire_5), .in(wire_6), .out(wire_39));
  TC_Switch # (.UUID(64'd1322051027298697595 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_12 (.en(wire_5), .in(wire_2), .out(wire_60));
  TC_Switch # (.UUID(64'd4279546958457643910 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_13 (.en(wire_5), .in(wire_52), .out(wire_8_0));
  TC_Switch # (.UUID(64'd1407183183188242545 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_14 (.en(wire_1), .in(wire_2), .out(wire_66));
  TC_Switch # (.UUID(64'd825188955478831971 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_15 (.en(wire_1), .in(wire_6), .out(wire_34));
  TC_Switch # (.UUID(64'd51925339328697175 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_16 (.en(wire_1), .in(wire_27), .out(wire_8_1));
  TC_Switch # (.UUID(64'd1175792227051955560 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_17 (.en(wire_4), .in(wire_6), .out(wire_37));
  TC_Switch # (.UUID(64'd1768630870230821680 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_18 (.en(wire_4), .in(wire_2), .out(wire_73));
  TC_Switch # (.UUID(64'd724522933239860619 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_19 (.en(wire_4), .in(wire_14), .out(wire_8_2));
  TC_Switch # (.UUID(64'd480414198129629098 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_20 (.en(wire_16), .in(wire_2), .out(wire_41));
  TC_Switch # (.UUID(64'd2236984552964180078 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_21 (.en(wire_16), .in(wire_6), .out(wire_71));
  TC_Switch # (.UUID(64'd2331894452996132707 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_16), .in(wire_36), .out(wire_8_3));
  TC_And # (.UUID(64'd4486090735793310582 ^ UUID), .BIT_WIDTH(64'd8)) And8_23 (.in0(wire_71), .in1(wire_41), .out(wire_36));
  TC_Nor # (.UUID(64'd428177551435513699 ^ UUID), .BIT_WIDTH(64'd8)) Nor8_24 (.in0(wire_37), .in1(wire_73), .out(wire_14));
  TC_Or # (.UUID(64'd1391410677810137682 ^ UUID), .BIT_WIDTH(64'd8)) Or8_25 (.in0(wire_39), .in1(wire_60), .out(wire_52));
  TC_Nand # (.UUID(64'd4025048423625330072 ^ UUID), .BIT_WIDTH(64'd8)) Nand8_26 (.in0(wire_34), .in1(wire_66), .out(wire_27));
  TC_Decoder3 # (.UUID(64'd3807680616509469728 ^ UUID)) Decoder3_27 (.dis(1'd0), .sel0(wire_69), .sel1(wire_42), .sel2(wire_31), .out0(wire_25), .out1(wire_30), .out2(wire_20), .out3(wire_75), .out4(wire_74), .out5(wire_46), .out6(wire_61), .out7(wire_70));
  TC_Xnor # (.UUID(64'd4268350311478768457 ^ UUID), .BIT_WIDTH(64'd8)) Xnor8_28 (.in0(wire_49), .in1(wire_81), .out(wire_59));
  TC_Xor # (.UUID(64'd4527214351160864442 ^ UUID), .BIT_WIDTH(64'd8)) Xor8_29 (.in0(wire_64), .in1(wire_12), .out(wire_40));
  TC_Not # (.UUID(64'd3618579806912338026 ^ UUID), .BIT_WIDTH(64'd8)) Not8_30 (.in(wire_58), .out(wire_63));
  TC_Mul # (.UUID(64'd86800450212264749 ^ UUID), .BIT_WIDTH(64'd8)) Mul8_31 (.in0(wire_51), .in1(wire_56), .out0(wire_80), .out1(wire_65));
  TC_Ashr # (.UUID(64'd4224934934216498493 ^ UUID), .BIT_WIDTH(64'd8)) Ashr8_32 (.in(wire_19), .shift(wire_53), .out(wire_43));
  TC_Neg # (.UUID(64'd687800544475925346 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_33 (.in(wire_11), .out(wire_67));
  TC_Rol # (.UUID(64'd1317775489477211882 ^ UUID), .BIT_WIDTH(64'd8)) Rol8_34 (.in(wire_47), .shift(wire_9), .out(wire_3));
  TC_Ror # (.UUID(64'd703554170280240747 ^ UUID), .BIT_WIDTH(64'd8)) Ror8_35 (.in(wire_76), .shift(wire_54), .out(wire_18));
  TC_Shr # (.UUID(64'd3748108855456900138 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_36 (.in(wire_17), .shift(wire_50), .out(wire_38));
  TC_Shl # (.UUID(64'd2176974598361832761 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_37 (.in(wire_85), .shift(wire_57), .out(wire_83));
  TC_Switch # (.UUID(64'd4483630066362025873 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_38 (.en(wire_0), .in(wire_2), .out(wire_12));
  TC_Switch # (.UUID(64'd3908274583674926227 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_39 (.en(wire_0), .in(wire_6), .out(wire_64));
  TC_Switch # (.UUID(64'd4553681126267151464 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_40 (.en(wire_0), .in(wire_40), .out(wire_8_5));
  TC_Switch # (.UUID(64'd4186982137889621636 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_41 (.en(wire_24), .in(wire_2), .out(wire_81));
  TC_Switch # (.UUID(64'd1386256187545231870 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_42 (.en(wire_24), .in(wire_6), .out(wire_49));
  TC_Switch # (.UUID(64'd2659168137376368183 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_43 (.en(wire_24), .in(wire_59), .out(wire_8_4));
  TC_Switch # (.UUID(64'd1704066470517955937 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_44 (.en(wire_26), .in(wire_6), .out(wire_58));
  TC_Switch # (.UUID(64'd2990116238052745508 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_45 (.en(wire_26), .in(wire_63), .out(wire_8_6));
  TC_Switch # (.UUID(64'd2820576902535906486 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_46 (.en(wire_5), .in(wire_2), .out(wire_53));
  TC_Switch # (.UUID(64'd59631099816967048 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_47 (.en(wire_5), .in(wire_6), .out(wire_19));
  TC_Switch # (.UUID(64'd3451848842388615139 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_5), .in(wire_43), .out(wire_22_3));
  TC_Switch # (.UUID(64'd4081918304701245721 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_49 (.en(wire_24), .in(wire_6), .out(wire_11));
  TC_Switch # (.UUID(64'd918819339348151073 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_50 (.en(wire_24), .in(wire_67), .out(wire_15_3));
  TC_Switch # (.UUID(64'd2919540118461118324 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_51 (.en(wire_1), .in(wire_6), .out(wire_79));
  TC_Switch # (.UUID(64'd3749247787192934141 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_52 (.en(wire_4), .in(wire_2), .out(wire_56));
  TC_Switch # (.UUID(64'd2395464300934186678 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_53 (.en(wire_4), .in(wire_6), .out(wire_51));
  TC_Switch # (.UUID(64'd1468357425860970596 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_54 (.en(wire_1), .in(wire_10), .out(wire_22_0));
  TC_Switch # (.UUID(64'd3788856213916320068 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_55 (.en(wire_1), .in(wire_78), .out(wire_44_0));
  TC_Switch # (.UUID(64'd3734865121253732914 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_56 (.en(wire_4), .in(wire_80), .out(wire_22_1));
  TC_Switch # (.UUID(64'd3847724417649658373 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_57 (.en(wire_4), .in(wire_65), .out(wire_44_1));
  TC_Switch # (.UUID(64'd2706629240204870554 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_58 (.en(wire_5), .in(wire_2), .out(wire_9));
  TC_Switch # (.UUID(64'd2001149239728006462 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_59 (.en(wire_5), .in(wire_6), .out(wire_47));
  TC_Switch # (.UUID(64'd2870113753177518410 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_60 (.en(wire_1), .in(wire_2), .out(wire_54));
  TC_Switch # (.UUID(64'd340004962580308093 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_61 (.en(wire_1), .in(wire_6), .out(wire_76));
  TC_Switch # (.UUID(64'd1684711578759063957 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_62 (.en(wire_4), .in(wire_6), .out(wire_17));
  TC_Switch # (.UUID(64'd2389968685784586327 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_63 (.en(wire_16), .in(wire_2), .out(wire_57));
  TC_Switch # (.UUID(64'd4535804765991235387 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_64 (.en(wire_16), .in(wire_6), .out(wire_85));
  TC_Switch # (.UUID(64'd667890680105453361 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_65 (.en(wire_4), .in(wire_2), .out(wire_50));
  TC_Switch # (.UUID(64'd3924371852208470488 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_66 (.en(wire_1), .in(wire_18), .out(wire_15_2));
  TC_Switch # (.UUID(64'd4550216520043673402 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_67 (.en(wire_5), .in(wire_3), .out(wire_15_4));
  TC_Switch # (.UUID(64'd1040267906917435020 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_68 (.en(wire_4), .in(wire_38), .out(wire_15_0));
  TC_Switch # (.UUID(64'd1068858050083309300 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_69 (.en(wire_16), .in(wire_83), .out(wire_15_1));
  TC_Switch # (.UUID(64'd1056292847970768806 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_70 (.en(wire_24), .in(wire_23), .out(wire_13_0));
  TC_Switch # (.UUID(64'd2775044829367273609 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_71 (.en(wire_16), .in(wire_21), .out(wire_13_1));
  TC_Switch # (.UUID(64'd683797453120618047 ^ UUID), .BIT_WIDTH(64'd8)) Output8z_72 (.en(wire_35), .in(wire_44), .out(D));
  TC_Switch # (.UUID(64'd1344327710761016922 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_73 (.en(wire_25), .in(wire_8), .out(wire_32_2));
  TC_Switch # (.UUID(64'd3164243025886628350 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_74 (.en(wire_30), .in(wire_22), .out(wire_32_1));
  TC_Switch # (.UUID(64'd389001382807605908 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_75 (.en(wire_20), .in(wire_15), .out(wire_32_0));
  TC_Or # (.UUID(64'd2298387723272408160 ^ UUID), .BIT_WIDTH(64'd1)) Or_76 (.in0(wire_1), .in1(wire_4), .out(wire_28));
  TC_And # (.UUID(64'd4016989336483643045 ^ UUID), .BIT_WIDTH(64'd1)) And_77 (.in0(wire_28), .in1(wire_30), .out(wire_35));
  TC_Mul # (.UUID(64'd3859724630390996553 ^ UUID), .BIT_WIDTH(64'd8)) DivMod8_78 (.in0(wire_79), .in1(wire_77), .out0(wire_10), .out1(wire_78));
  TC_Switch # (.UUID(64'd2129354784258529228 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_79 (.en(wire_1), .in(wire_2), .out());
  TC_Constant # (.UUID(64'd1325873776756270234 ^ UUID), .BIT_WIDTH(64'd8), .value(8'hAA)) Constant8_80 (.out(wire_77));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [7:0] wire_2;
  assign wire_2 = B;
  wire [7:0] wire_3;
  wire [0:0] wire_4;
  wire [0:0] wire_5;
  wire [7:0] wire_6;
  assign wire_6 = A;
  wire [0:0] wire_7;
  wire [7:0] wire_8;
  wire [7:0] wire_8_0;
  wire [7:0] wire_8_1;
  wire [7:0] wire_8_2;
  wire [7:0] wire_8_3;
  wire [7:0] wire_8_4;
  wire [7:0] wire_8_5;
  wire [7:0] wire_8_6;
  assign wire_8 = wire_8_0|wire_8_1|wire_8_2|wire_8_3|wire_8_4|wire_8_5|wire_8_6;
  wire [7:0] wire_9;
  wire [7:0] wire_10;
  wire [7:0] wire_11;
  wire [7:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_13_0;
  wire [0:0] wire_13_1;
  assign wire_13 = wire_13_0|wire_13_1;
  assign CF = wire_13;
  wire [7:0] wire_14;
  wire [7:0] wire_15;
  wire [7:0] wire_15_0;
  wire [7:0] wire_15_1;
  wire [7:0] wire_15_2;
  wire [7:0] wire_15_3;
  wire [7:0] wire_15_4;
  assign wire_15 = wire_15_0|wire_15_1|wire_15_2|wire_15_3|wire_15_4;
  wire [0:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_18;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  wire [7:0] wire_22_0;
  wire [7:0] wire_22_1;
  wire [7:0] wire_22_2;
  wire [7:0] wire_22_3;
  wire [7:0] wire_22_4;
  assign wire_22 = wire_22_0|wire_22_1|wire_22_2|wire_22_3|wire_22_4;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [7:0] wire_27;
  wire [0:0] wire_28;
  wire [7:0] wire_29;
  assign wire_29 = Instruction;
  wire [0:0] wire_30;
  wire [0:0] wire_31;
  wire [7:0] wire_32;
  wire [7:0] wire_32_0;
  wire [7:0] wire_32_1;
  wire [7:0] wire_32_2;
  assign wire_32 = wire_32_0|wire_32_1|wire_32_2;
  assign C = wire_32;
  wire [7:0] wire_33;
  wire [7:0] wire_34;
  wire [0:0] wire_35;
  assign D_OUT_EN = wire_35;
  wire [7:0] wire_36;
  wire [7:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [7:0] wire_40;
  wire [7:0] wire_41;
  wire [0:0] wire_42;
  wire [7:0] wire_43;
  wire [7:0] wire_44;
  wire [7:0] wire_44_0;
  wire [7:0] wire_44_1;
  assign wire_44 = wire_44_0|wire_44_1;
  wire [7:0] wire_45;
  wire [0:0] wire_46;
  wire [7:0] wire_47;
  wire [0:0] wire_48;
  wire [7:0] wire_49;
  wire [7:0] wire_50;
  wire [7:0] wire_51;
  wire [7:0] wire_52;
  wire [7:0] wire_53;
  wire [7:0] wire_54;
  wire [0:0] wire_55;
  wire [7:0] wire_56;
  wire [7:0] wire_57;
  wire [7:0] wire_58;
  wire [7:0] wire_59;
  wire [7:0] wire_60;
  wire [0:0] wire_61;
  wire [7:0] wire_62;
  wire [7:0] wire_63;
  wire [7:0] wire_64;
  wire [7:0] wire_65;
  wire [7:0] wire_66;
  wire [7:0] wire_67;
  wire [7:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [7:0] wire_71;
  wire [7:0] wire_72;
  wire [7:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [7:0] wire_76;
  wire [7:0] wire_77;
  wire [7:0] wire_78;
  wire [7:0] wire_79;
  wire [7:0] wire_80;
  wire [7:0] wire_81;
  wire [0:0] wire_82;
  wire [7:0] wire_83;
  wire [7:0] wire_84;
  wire [7:0] wire_85;
  wire [7:0] wire_86;

endmodule
