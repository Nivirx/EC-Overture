module ECP8e (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_Switch # (.UUID(64'd1715727152826423794 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_0 (.en(wire_50), .in(wire_48), .out(wire_41));
  TC_Halt # (.UUID(64'd2976448359382631736 ^ UUID)) Halt_1 (.clk(clk), .rst(rst), .en(wire_67));
  TC_Not # (.UUID(64'd2472047754744094114 ^ UUID), .BIT_WIDTH(64'd1)) Not_2 (.in(wire_61), .out(wire_67));
  TC_IOSwitch # (.UUID(64'd2352853726822514667 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_3 (.in(wire_56), .en(wire_38), .out(arch_output_value));
  TC_Program8_1 # (.UUID(64'd2319742357034652024 ^ UUID), .DEFAULT_FILE_NAME("outport_test.bin"), .ARG_SIG("outport_test=%s")) Program8_1_4 (.clk(clk), .rst(rst), .address(wire_5), .out(wire_48));
  TC_Switch # (.UUID(64'd556654018140205888 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_5 (.en(wire_27), .in(arch_input_value), .out(wire_39));
  ALU # (.UUID(64'd3424272698184478142 ^ UUID)) ALU_6 (.clk(clk), .rst(rst), .Instruction(wire_41), .A(wire_35), .B(wire_75), .D_OUT_EN(wire_15), .D(wire_71), .CF(), .C(wire_66));
  TC_Ram # (.UUID(64'd1661974221341126710 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd64)) Ram_7 (.clk(clk), .rst(rst), .load(1'd0), .save(1'd0), .address(32'd0), .in0(64'd0), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(), .out1(), .out2(), .out3());
  TC_Buffer # (.UUID(64'd3602924629092547678 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_8 (.in(wire_48), .out(wire_28));
  TC_Buffer # (.UUID(64'd1036402492479265627 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_9 (.in(wire_1), .out(wire_55));
  TC_Buffer # (.UUID(64'd3234323155509956945 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_10 (.in(wire_23), .out(wire_60));
  TC_Buffer # (.UUID(64'd2118082778336995084 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_11 (.in(wire_18), .out(wire_77));
  TC_Buffer # (.UUID(64'd3247628008814229228 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_12 (.in(wire_20), .out(wire_72));
  TC_Buffer # (.UUID(64'd3783645420539942969 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_13 (.in(wire_33), .out(wire_73));
  TC_Buffer # (.UUID(64'd101493406757515111 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_14 (.in(wire_31), .out(wire_43));
  TC_Buffer # (.UUID(64'd1648258134768700275 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_15 (.in(wire_2), .out(wire_56));
  TC_Buffer # (.UUID(64'd297196408869131089 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_16 (.in(wire_39), .out(wire_51));
  TC_Decoder3 # (.UUID(64'd319890292667874856 ^ UUID)) Decoder3_17 (.dis(wire_19), .sel0(wire_47), .sel1(wire_69), .sel2(wire_70), .out0(wire_32), .out1(wire_34), .out2(wire_46), .out3(wire_9), .out4(wire_7), .out5(wire_62), .out6(wire_26), .out7(wire_53));
  TC_Decoder3 # (.UUID(64'd4421418411989485663 ^ UUID)) Decoder3_18 (.dis(wire_19), .sel0(wire_52), .sel1(wire_58), .sel2(wire_4), .out0(wire_65), .out1(wire_44), .out2(wire_59), .out3(wire_54), .out4(wire_14), .out5(wire_21), .out6(wire_24), .out7(wire_42));
  TC_Splitter8 # (.UUID(64'd274394922392375603 ^ UUID)) Splitter8_19 (.in(wire_28), .out0(wire_52), .out1(wire_58), .out2(wire_4), .out3(wire_47), .out4(wire_69), .out5(wire_70), .out6(), .out7());
  TC_Maker16 # (.UUID(64'd4271331395148101399 ^ UUID)) Maker16_20 (.in0(wire_23), .in1(wire_18), .out(wire_64));
  TC_Xor # (.UUID(64'd4015117391550831776 ^ UUID), .BIT_WIDTH(64'd1)) Xor_21 (.in0(wire_45), .in1(wire_65), .out(wire_68));
  TC_Switch # (.UUID(64'd4445417212749692549 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_22 (.en(wire_26), .in(wire_51), .out(wire_6_1));
  TC_Switch # (.UUID(64'd556730729123347464 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_23 (.en(wire_24), .in(wire_17), .out(wire_2));
  TC_Buffer # (.UUID(64'd3347726601253752187 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_24 (.in(wire_10), .out(wire_50));
  TC_Switch # (.UUID(64'd1860343635038049181 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_25 (.en(wire_8), .in(wire_17), .out(wire_6_0));
  TC_Or # (.UUID(64'd4336129294321593228 ^ UUID), .BIT_WIDTH(64'd1)) Or_26 (.in0(wire_25), .in1(wire_3), .out(wire_45));
  TC_Xor # (.UUID(64'd1518074666294394017 ^ UUID), .BIT_WIDTH(64'd1)) Xor_27 (.in0(wire_54), .in1(wire_10), .out(wire_12));
  TC_Nand # (.UUID(64'd3859693831101792233 ^ UUID), .BIT_WIDTH(64'd1)) Nand_28 (.in0(wire_42), .in1(wire_53), .out(wire_22));
  TC_Switch # (.UUID(64'd1247979186234576792 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_29 (.en(wire_3), .in(wire_28), .out(wire_6_4));
  TC_Or3 # (.UUID(64'd4011049292989256787 ^ UUID), .BIT_WIDTH(64'd1)) Or3_30 (.in0(wire_3), .in1(wire_10), .in2(wire_25), .out(wire_19));
  TC_Switch # (.UUID(64'd2893193334261668714 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_31 (.en(wire_10), .in(wire_16), .out(wire_6_3));
  TC_And # (.UUID(64'd3005434726623612484 ^ UUID), .BIT_WIDTH(64'd1)) And_32 (.in0(wire_25), .in1(wire_76), .out(wire_49));
  TC_Switch # (.UUID(64'd929078426947889085 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_33 (.en(wire_25), .in(wire_28), .out(wire_63));
  TC_Counter # (.UUID(64'd3263272588803768522 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_34 (.clk(clk), .rst(rst), .save(wire_49), .in(wire_1), .out(wire_5));
  TC_Buffer # (.UUID(64'd2235373354836046298 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_35 (.in(wire_22), .out(wire_61));
  TC_Buffer # (.UUID(64'd2032593801523540386 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_36 (.in(wire_5), .out());
  TC_Buffer # (.UUID(64'd2286316240340576623 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_37 (.in(wire_15), .out(wire_36));
  TC_Splitter16 # (.UUID(64'd2817158020377327923 ^ UUID)) Splitter16_38 (.in(wire_29), .out0(wire_16), .out1(wire_0));
  TC_Switch # (.UUID(64'd2251356442933710957 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_39 (.en(wire_36), .in(wire_0), .out(wire_6_2));
  TC_Buffer # (.UUID(64'd2774123988237700806 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_40 (.in(wire_24), .out(wire_38));
  TC_Buffer # (.UUID(64'd2259435457617166464 ^ UUID), .BIT_WIDTH(64'd1)) Buffer1_41 (.in(wire_26), .out(wire_27));
  TC_Nor # (.UUID(64'd28166036220749041 ^ UUID), .BIT_WIDTH(64'd1)) Nor_42 (.in0(wire_26), .in1(wire_24), .out(wire_37));
  TC_And # (.UUID(64'd2711603589399634934 ^ UUID), .BIT_WIDTH(64'd1)) And_43 (.in0(wire_40), .in1(wire_37), .out(wire_8));
  TC_Splitter16 # (.UUID(64'd4364533521657012903 ^ UUID)) Splitter16_44 (.in(wire_74), .out0(wire_11), .out1(wire_30));
  TC_Buffer # (.UUID(64'd1306800471778976915 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_45 (.in(wire_11), .out(wire_35));
  TC_Buffer # (.UUID(64'd4600618263124473635 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_46 (.in(wire_30), .out(wire_75));
  TC_Switch # (.UUID(64'd2102499097582599256 ^ UUID), .BIT_WIDTH(64'd16)) Switch16_47 (.en(wire_10), .in(wire_64), .out(wire_74));
  TC_Buffer # (.UUID(64'd1794452372346720268 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_48 (.in(wire_66), .out(wire_57));
  TC_Buffer # (.UUID(64'd3772267359649597453 ^ UUID), .BIT_WIDTH(64'd8)) Buffer8_49 (.in(wire_71), .out(wire_13));
  TC_Maker16 # (.UUID(64'd1181495850574424 ^ UUID)) Maker16_50 (.in0(wire_57), .in1(wire_13), .out(wire_29));
  RegisterPlus # (.UUID(64'd2661760033600874299 ^ UUID)) RegisterPlus_51 (.clk(clk), .rst(rst), .Load(wire_32), .Save_value(wire_6), .Save(wire_68), .Always_output(wire_1), .Output(wire_17_4));
  RegisterPlus # (.UUID(64'd2163217265803647012 ^ UUID)) RegisterPlus_52 (.clk(clk), .rst(rst), .Load(wire_34), .Save_value(wire_6), .Save(wire_44), .Always_output(wire_23), .Output(wire_17_5));
  RegisterPlus # (.UUID(64'd1347627285814452637 ^ UUID)) RegisterPlus_53 (.clk(clk), .rst(rst), .Load(wire_46), .Save_value(wire_6), .Save(wire_59), .Always_output(wire_18), .Output(wire_17_3));
  RegisterPlus # (.UUID(64'd3166915688793493761 ^ UUID)) RegisterPlus_54 (.clk(clk), .rst(rst), .Load(wire_9), .Save_value(wire_6), .Save(wire_12), .Always_output(wire_20), .Output(wire_17_2));
  RegisterPlus # (.UUID(64'd4519434156825869138 ^ UUID)) RegisterPlus_55 (.clk(clk), .rst(rst), .Load(wire_7), .Save_value(wire_6), .Save(wire_14), .Always_output(wire_33), .Output(wire_17_1));
  RegisterPlus # (.UUID(64'd3857793667730710479 ^ UUID)) RegisterPlus_56 (.clk(clk), .rst(rst), .Load(wire_62), .Save_value(wire_6), .Save(wire_21), .Always_output(wire_31), .Output(wire_17_0));
  DEC # (.UUID(64'd3963022757837899629 ^ UUID)) DEC_57 (.clk(clk), .rst(rst), .Instruction(wire_28), .IMM_EN(wire_3), .ALU_EN(wire_10), .COPY_EN(wire_40), .BRANCH_EN(wire_25));
  COND # (.UUID(64'd1986738645304097046 ^ UUID)) COND_58 (.clk(clk), .rst(rst), .Condition(wire_63), .Input(wire_20), .Result(wire_76));

  wire [7:0] wire_0;
  wire [7:0] wire_1;
  wire [7:0] wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_6;
  wire [7:0] wire_6_0;
  wire [7:0] wire_6_1;
  wire [7:0] wire_6_2;
  wire [7:0] wire_6_3;
  wire [7:0] wire_6_4;
  assign wire_6 = wire_6_0|wire_6_1|wire_6_2|wire_6_3|wire_6_4;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [7:0] wire_11;
  wire [0:0] wire_12;
  wire [7:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_17_0;
  wire [7:0] wire_17_1;
  wire [7:0] wire_17_2;
  wire [7:0] wire_17_3;
  wire [7:0] wire_17_4;
  wire [7:0] wire_17_5;
  assign wire_17 = wire_17_0|wire_17_1|wire_17_2|wire_17_3|wire_17_4|wire_17_5;
  wire [7:0] wire_18;
  wire [0:0] wire_19;
  wire [7:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [7:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  assign arch_input_enable = wire_27;
  wire [7:0] wire_28;
  wire [15:0] wire_29;
  wire [7:0] wire_30;
  wire [7:0] wire_31;
  wire [0:0] wire_32;
  wire [7:0] wire_33;
  wire [0:0] wire_34;
  wire [7:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  assign arch_output_enable = wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [7:0] wire_41;
  wire [0:0] wire_42;
  wire [7:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [7:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [7:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [7:0] wire_55;
  wire [7:0] wire_56;
  wire [7:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [7:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [7:0] wire_63;
  wire [15:0] wire_64;
  wire [0:0] wire_65;
  wire [7:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [7:0] wire_71;
  wire [7:0] wire_72;
  wire [7:0] wire_73;
  wire [15:0] wire_74;
  wire [7:0] wire_75;
  wire [0:0] wire_76;
  wire [7:0] wire_77;

endmodule
